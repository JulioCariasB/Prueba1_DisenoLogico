// VGA protocol constants for 640x480 resolution
`define VGA_WIDTH  640
`define VGA_HEIGHT 480
`define VGA_HLIMIT 800
`define VGA_VLIMIT 525
`define VGA_HSYNC_PULSE_START 656
`define VGA_HSYNC_PULSE_END   752
`define VGA_VSYNC_PULSE_START 490
`define VGA_VSYNC_PULSE_END   492

`define COLOR_BITS 8
