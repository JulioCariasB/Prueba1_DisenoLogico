/*
TODO: Instantiate VGA640x480 module 
TODO: Instantiate VGAClock module 
TODO: Connect the two modules 
*/
